`include "vutils_macros.svh"

// verif utils package
package vutils_pkg;
  `include "vutils_types.svh"
endpackage // vutils_pkg
